module Ins_mem (
    input [31:0] adr,
    output reg [31:0] dout
);

wire [4:0] cmd = adr[4:0];
always@(*) begin
        case(cmd)
        
        4'b0000: dout = 32'b101000_01001_01001_0000000000000000;
        4'b0001: dout = 32'b101000_01010_01010_0000000000000001;
        4'b0010: dout = 32'b101000_01011_01011_0000000000000000;
        4'b0011: dout = 32'b101000_01100_01100_0000000000010100;
        4'b0100: dout = 32'b000000_01001_01010_10001_00000_100000;
        4'b0101: dout = 32'b101000_01001_01010_0000000000000000;
        4'b0110: dout = 32'b101000_01010_10001_0000000000000000;
        4'b0111: dout = 32'b101000_01011_01011_0000000000000010;
        4'b1000: dout = 32'b000100_01100_01011_0000000000000110;
        4'b1001: dout = 32'b100110_00000000000000000000000101;
        4'b1010: dout = 32'b101011_01100_10001_0000000000000101;
        4'b1011: dout = 32'b000000_01100_10001_10010_00000_101010;
        
        default : dout =32'dx;
        endcase
    end
    
endmodule
